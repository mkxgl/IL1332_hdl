`timescale 1ns / 1ps
module nand2_delay(
	input logic a,
	input logic b,
	output logic y
	);

	assign #1ns y = ~(a&b);

endmodule